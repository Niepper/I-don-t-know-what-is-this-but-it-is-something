module main


fn main() {
	animal := ["wild dog", "wolf", "gryphon", "Strzyga", "dragon", "devil"]

	println(animal[(167-1)%6])
}
